//
// Acquire data from one ADC 3424
//
// Four channels -> four ADC waveforms, four discriminators
//

module adc_discr_group
 (
  input[7:0] adc_DP,
  input[7:0] adc_DM,
 );

 endmodule
